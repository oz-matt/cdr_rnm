`ifndef NREAL_GUARD
`define NREAL_GUARD

package nreal;

  nettype real nreal;

endpackage

`endif
