
`include "top_test.sv"

