`ifndef EENET_SYMBOLS_GUARD
`define EENET_SYMBOLS_GUARD

`include "VsrcG.sv"
`include "VRsrc.sv"
`include "Isrc.sv"
`include "IsrcG.sv"
`include "ResG.sv"
`include "CapG.sv"
`endif
